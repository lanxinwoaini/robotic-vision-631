-------------------------------------------------------------------------------
-- Inverse ROMs
--
-- DESCRIPTION
--
-- Two ROMs containing 1/1 .. 1/255 in 8.16 fixed point
-- (6kb � 384 LUTs each, 128 CLBs)
--
-- VERSION SPECIFIC INFORMATION
--
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;
--use ieee.std_logic_signed.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following lines to use the declarations that are
-- provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity inv_table is
port (
value_A : in std_logic_vector(7 downto 0);
value_B : in std_logic_vector(7 downto 0);
inverse_A : out std_logic_vector(23 downto 0);
inverse_B : out std_logic_vector(23 downto 0)
);
end inv_table;

architecture Behavioral of inv_table is
	subtype inverse_word is std_logic_vector(23 downto 0);
	type inverse_table is array (0 to 255) of inverse_word;
	constant inverses : inverse_table := inverse_table'(
		inverse_word'("000000000000000000000000"),
		inverse_word'("000011111111000000000000"),
		inverse_word'("000001111111100000000000"),
		inverse_word'("000001010101000000000000"),
		inverse_word'("000000111111110000000000"),
		inverse_word'("000000110011000000000000"),
		inverse_word'("000000101010100000000000"),
		inverse_word'("000000100100011011011011"),
		inverse_word'("000000011111111000000000"),
		inverse_word'("000000011100010101010101"),
		inverse_word'("000000011001100000000000"),
		inverse_word'("000000010111001011101001"),
		inverse_word'("000000010101010000000000"),
		inverse_word'("000000010011100111011001"),
		inverse_word'("000000010010001101101110"),
		inverse_word'("000000010001000000000000"),
		inverse_word'("000000001111111100000000"),
		inverse_word'("000000001111000000000000"),
		inverse_word'("000000001110001010101011"),
		inverse_word'("000000001101011010111101"),
		inverse_word'("000000001100110000000000"),
		inverse_word'("000000001100001001001001"),
		inverse_word'("000000001011100101110100"),
		inverse_word'("000000001011000101100100"),
		inverse_word'("000000001010101000000000"),
		inverse_word'("000000001010001100110011"),
		inverse_word'("000000001001110011101100"),
		inverse_word'("000000001001011100011100"),
		inverse_word'("000000001001000110110111"),
		inverse_word'("000000001000110010110001"),
		inverse_word'("000000001000100000000000"),
		inverse_word'("000000001000001110011101"),
		inverse_word'("000000000111111110000000"),
		inverse_word'("000000000111101110100011"),
		inverse_word'("000000000111100000000000"),
		inverse_word'("000000000111010010010010"),
		inverse_word'("000000000111000101010101"),
		inverse_word'("000000000110111001000101"),
		inverse_word'("000000000110101101011110"),
		inverse_word'("000000000110100010011110"),
		inverse_word'("000000000110011000000000"),
		inverse_word'("000000000110001110000011"),
		inverse_word'("000000000110000100100101"),
		inverse_word'("000000000101111011100010"),
		inverse_word'("000000000101110010111010"),
		inverse_word'("000000000101101010101011"),
		inverse_word'("000000000101100010110010"),
		inverse_word'("000000000101011011001111"),
		inverse_word'("000000000101010100000000"),
		inverse_word'("000000000101001101000100"),
		inverse_word'("000000000101000110011010"),
		inverse_word'("000000000101000000000000"),
		inverse_word'("000000000100111001110110"),
		inverse_word'("000000000100110011111011"),
		inverse_word'("000000000100101110001110"),
		inverse_word'("000000000100101000101111"),
		inverse_word'("000000000100100011011011"),
		inverse_word'("000000000100011110010100"),
		inverse_word'("000000000100011001011000"),
		inverse_word'("000000000100010100100111"),
		inverse_word'("000000000100010000000000"),
		inverse_word'("000000000100001011100011"),
		inverse_word'("000000000100000111001110"),
		inverse_word'("000000000100000011000011"),
		inverse_word'("000000000011111111000000"),
		inverse_word'("000000000011111011000101"),
		inverse_word'("000000000011110111010001"),
		inverse_word'("000000000011110011100101"),
		inverse_word'("000000000011110000000000"),
		inverse_word'("000000000011101100100001"),
		inverse_word'("000000000011101001001001"),
		inverse_word'("000000000011100101110111"),
		inverse_word'("000000000011100010101011"),
		inverse_word'("000000000011011111100100"),
		inverse_word'("000000000011011100100011"),
		inverse_word'("000000000011011001100110"),
		inverse_word'("000000000011010110101111"),
		inverse_word'("000000000011010011111101"),
		inverse_word'("000000000011010001001111"),
		inverse_word'("000000000011001110100101"),
		inverse_word'("000000000011001100000000"),
		inverse_word'("000000000011001001011111"),
		inverse_word'("000000000011000111000010"),
		inverse_word'("000000000011000100101000"),
		inverse_word'("000000000011000010010010"),
		inverse_word'("000000000011000000000000"),
		inverse_word'("000000000010111101110001"),
		inverse_word'("000000000010111011100110"),
		inverse_word'("000000000010111001011101"),
		inverse_word'("000000000010110111011000"),
		inverse_word'("000000000010110101010101"),
		inverse_word'("000000000010110011010110"),
		inverse_word'("000000000010110001011001"),
		inverse_word'("000000000010101111011111"),
		inverse_word'("000000000010101101100111"),
		inverse_word'("000000000010101011110011"),
		inverse_word'("000000000010101010000000"),
		inverse_word'("000000000010101000010000"),
		inverse_word'("000000000010100110100010"),
		inverse_word'("000000000010100100110110"),
		inverse_word'("000000000010100011001101"),
		inverse_word'("000000000010100001100101"),
		inverse_word'("000000000010100000000000"),
		inverse_word'("000000000010011110011101"),
		inverse_word'("000000000010011100111011"),
		inverse_word'("000000000010011011011011"),
		inverse_word'("000000000010011001111110"),
		inverse_word'("000000000010011000100001"),
		inverse_word'("000000000010010111000111"),
		inverse_word'("000000000010010101101110"),
		inverse_word'("000000000010010100010111"),
		inverse_word'("000000000010010011000010"),
		inverse_word'("000000000010010001101110"),
		inverse_word'("000000000010010000011011"),
		inverse_word'("000000000010001111001010"),
		inverse_word'("000000000010001101111010"),
		inverse_word'("000000000010001100101100"),
		inverse_word'("000000000010001011011111"),
		inverse_word'("000000000010001010010100"),
		inverse_word'("000000000010001001001001"),
		inverse_word'("000000000010001000000000"),
		inverse_word'("000000000010000110111000"),
		inverse_word'("000000000010000101110001"),
		inverse_word'("000000000010000100101100"),
		inverse_word'("000000000010000011100111"),
		inverse_word'("000000000010000010100100"),
		inverse_word'("000000000010000001100010"),
		inverse_word'("000000000010000000100000"),
		inverse_word'("000000000001111111100000"),
		inverse_word'("000000000001111110100001"),
		inverse_word'("000000000001111101100010"),
		inverse_word'("000000000001111100100101"),
		inverse_word'("000000000001111011101001"),
		inverse_word'("000000000001111010101101"),
		inverse_word'("000000000001111001110011"),
		inverse_word'("000000000001111000111001"),
		inverse_word'("000000000001111000000000"),
		inverse_word'("000000000001110111001000"),
		inverse_word'("000000000001110110010001"),
		inverse_word'("000000000001110101011010"),
		inverse_word'("000000000001110100100101"),
		inverse_word'("000000000001110011110000"),
		inverse_word'("000000000001110010111011"),
		inverse_word'("000000000001110010001000"),
		inverse_word'("000000000001110001010101"),
		inverse_word'("000000000001110000100011"),
		inverse_word'("000000000001101111110010"),
		inverse_word'("000000000001101111000001"),
		inverse_word'("000000000001101110010001"),
		inverse_word'("000000000001101101100010"),
		inverse_word'("000000000001101100110011"),
		inverse_word'("000000000001101100000101"),
		inverse_word'("000000000001101011011000"),
		inverse_word'("000000000001101010101011"),
		inverse_word'("000000000001101001111110"),
		inverse_word'("000000000001101001010011"),
		inverse_word'("000000000001101000100111"),
		inverse_word'("000000000001100111111101"),
		inverse_word'("000000000001100111010011"),
		inverse_word'("000000000001100110101001"),
		inverse_word'("000000000001100110000000"),
		inverse_word'("000000000001100101010111"),
		inverse_word'("000000000001100100101111"),
		inverse_word'("000000000001100100001000"),
		inverse_word'("000000000001100011100001"),
		inverse_word'("000000000001100010111010"),
		inverse_word'("000000000001100010010100"),
		inverse_word'("000000000001100001101110"),
		inverse_word'("000000000001100001001001"),
		inverse_word'("000000000001100000100100"),
		inverse_word'("000000000001100000000000"),
		inverse_word'("000000000001011111011100"),
		inverse_word'("000000000001011110111001"),
		inverse_word'("000000000001011110010101"),
		inverse_word'("000000000001011101110011"),
		inverse_word'("000000000001011101010000"),
		inverse_word'("000000000001011100101111"),
		inverse_word'("000000000001011100001101"),
		inverse_word'("000000000001011011101100"),
		inverse_word'("000000000001011011001011"),
		inverse_word'("000000000001011010101011"),
		inverse_word'("000000000001011010001011"),
		inverse_word'("000000000001011001101011"),
		inverse_word'("000000000001011001001100"),
		inverse_word'("000000000001011000101101"),
		inverse_word'("000000000001011000001110"),
		inverse_word'("000000000001010111101111"),
		inverse_word'("000000000001010111010001"),
		inverse_word'("000000000001010110110100"),
		inverse_word'("000000000001010110010110"),
		inverse_word'("000000000001010101111001"),
		inverse_word'("000000000001010101011100"),
		inverse_word'("000000000001010101000000"),
		inverse_word'("000000000001010100100100"),
		inverse_word'("000000000001010100001000"),
		inverse_word'("000000000001010011101100"),
		inverse_word'("000000000001010011010001"),
		inverse_word'("000000000001010010110110"),
		inverse_word'("000000000001010010011011"),
		inverse_word'("000000000001010010000001"),
		inverse_word'("000000000001010001100110"),
		inverse_word'("000000000001010001001100"),
		inverse_word'("000000000001010000110011"),
		inverse_word'("000000000001010000011001"),
		inverse_word'("000000000001010000000000"),
		inverse_word'("000000000001001111100111"),
		inverse_word'("000000000001001111001110"),
		inverse_word'("000000000001001110110110"),
		inverse_word'("000000000001001110011110"),
		inverse_word'("000000000001001110000110"),
		inverse_word'("000000000001001101101110"),
		inverse_word'("000000000001001101010110"),
		inverse_word'("000000000001001100111111"),
		inverse_word'("000000000001001100101000"),
		inverse_word'("000000000001001100010001"),
		inverse_word'("000000000001001011111010"),
		inverse_word'("000000000001001011100100"),
		inverse_word'("000000000001001011001101"),
		inverse_word'("000000000001001010110111"),
		inverse_word'("000000000001001010100001"),
		inverse_word'("000000000001001010001100"),
		inverse_word'("000000000001001001110110"),
		inverse_word'("000000000001001001100001"),
		inverse_word'("000000000001001001001100"),
		inverse_word'("000000000001001000110111"),
		inverse_word'("000000000001001000100010"),
		inverse_word'("000000000001001000001110"),
		inverse_word'("000000000001000111111001"),
		inverse_word'("000000000001000111100101"),
		inverse_word'("000000000001000111010001"),
		inverse_word'("000000000001000110111101"),
		inverse_word'("000000000001000110101010"),
		inverse_word'("000000000001000110010110"),
		inverse_word'("000000000001000110000011"),
		inverse_word'("000000000001000101110000"),
		inverse_word'("000000000001000101011101"),
		inverse_word'("000000000001000101001010"),
		inverse_word'("000000000001000100110111"),
		inverse_word'("000000000001000100100101"),
		inverse_word'("000000000001000100010010"),
		inverse_word'("000000000001000100000000"),
		inverse_word'("000000000001000011101110"),
		inverse_word'("000000000001000011011100"),
		inverse_word'("000000000001000011001010"),
		inverse_word'("000000000001000010111001"),
		inverse_word'("000000000001000010100111"),
		inverse_word'("000000000001000010010110"),
		inverse_word'("000000000001000010000101"),
		inverse_word'("000000000001000001110100"),
		inverse_word'("000000000001000001100011"),
		inverse_word'("000000000001000001010010"),
		inverse_word'("000000000001000001000001"),
		inverse_word'("000000000001000000110001"),
		inverse_word'("000000000001000000100000"),
		inverse_word'("000000000001000000010000"),
		inverse_word'("000000000001000000000000"));
begin
	inverse_A <= inverses(conv_integer("0" &  value_A));
	inverse_B <= inverses(conv_integer("0" &  value_B));
end Behavioral;